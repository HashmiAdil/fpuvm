// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: types_bus0 
package sv_types_bus0; 
  parameter CFG_BUS0_XSLV_BOOTROM = 0;
  parameter CFG_BUS0_XSLV_ROMIMAGE = 1;
  parameter CFG_BUS0_XSLV_SRAM = 2;
  parameter CFG_BUS0_XSLV_UART1 = 3;
  parameter CFG_BUS0_XSLV_GPIO = 4;
  parameter CFG_BUS0_XSLV_IRQCTRL = 5;
  parameter CFG_BUS0_XSLV_GNSS_SS = 6;
  parameter CFG_BUS0_XSLV_EXTFLASH = 7;
  parameter CFG_BUS0_XSLV_ETHMAC = 8;
  parameter CFG_BUS0_XSLV_DSU = 9;
  parameter CFG_BUS0_XSLV_GPTIMERS = 10;
  parameter CFG_BUS0_XSLV_OTP = 11;
  parameter CFG_BUS0_XSLV_PNP = 12;
  parameter CFG_BUS0_XSLV_TOTAL = 13;
  parameter CFG_BUS0_XMST_WORKGROUP = 0;
  parameter CFG_BUS0_XMST_ETHMAC = 1;
  parameter CFG_BUS0_XMST_MSTUART = 2;
  parameter CFG_BUS0_XMST_DMI = 3;
  parameter CFG_BUS0_XMST_TOTAL = 4;
endpackage : sv_types_bus0 

import sv_types_bus0::* 

