// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: types_misc 
package sv_types_misc; 
  parameter CFG_IRQ_UNUSED = 0;
  parameter CFG_IRQ_UART1 = 1;
  parameter CFG_IRQ_ETHMAC = 2;
  parameter CFG_IRQ_GPTIMERS = 3;
  parameter CFG_IRQ_GNSSENGINE = 4;
  parameter CFG_IRQ_TOTAL = 5;
  parameter spi_out_none = 5;
endpackage : sv_types_misc 

import sv_types_misc::* 

